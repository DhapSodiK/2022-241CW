// Task 3 - 2022
module task3;

#(output logic [8:0] Q, input logic CLK, n_RESET, DATAIN);

always_ff @(posedge CLK)	begin
if (counter == 0) begin

end

endmodule
